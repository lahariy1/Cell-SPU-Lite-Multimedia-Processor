package definitions;
	parameter WORD = 32;
	parameter HALF_WORD = 16;
	parameter BYTE = 8;
	parameter QUAD_WORD = 128;
	parameter NIBBLE = 4;
	
	parameter SMAX = $bitstoshortreal(32'h7fffffff);
	parameter SMIN = $bitstoshortreal(32'h80000000);
	
	parameter EVEN = 0;
	parameter ODD = 1;
	
	typedef enum logic[10:0] {
							ADD_HALFWORD 			 	 					= 11'b00011001000,
							ADD_HALFWORD_IMMEDIATE   	 					= 11'b00011101000,
							ADD_WORD				  						= 11'b00011000000,
							ADD_WORD_IMMEDIATE        						= 11'b00011100000,
							SUB_FROM_HALFWORD		 						= 11'b00001001000,
							SUB_FROM_HALFWORD_IMMEDIATE						= 11'b00001101000,
							SUB_FROM_WORD			 						= 11'b00001000000,
							SUB_FROM_WORD_IMMEDIATE							= 11'b00001100000,
							MULTIPLY 				  						= 11'b01111000100,
							MULITPLY_UNSIGNED		  						= 11'b01111001100,
							MULTIPLY_IMMEDIATE		  						= 11'b01110100000,
							MULTIPLY_AND_ADD		  						= 11'b11000000000,
							COUNTING_LEADING_ZEROS	  						= 11'b01010100101,
							FORM_SELECT_MASK_BYTES_IMMEDIATE				= 11'b00110010100,
							FORM_SELECT_MASK_BYTES   						= 11'b00110110110,
							FORM_SELECT_MASK_HALFWORD 						= 11'b00110110101,
							FORM_SELECT_MASK_WORD	 						= 11'b00110110100,
							AND						  						= 11'b00011000001,
							AND_HALFWORD_IMMEDIATE	  						= 11'b00010101000,
							AND_WORD_IMMEDIATE		  						= 11'b00010100000,
							OR					  							= 11'b00001000001,
							OR_BYTE_IMMEDIATE								= 11'b00000110000,
							OR_HALFWORD_IMMEDIATE	  						= 11'b00000101000,
							OR_WORD_IMMEDIATE	      						= 11'b00000100000,
							NOR						  						= 11'b00001001001,
							XOR						  						= 11'b01001000001,
							XOR_BYTE_IMMEDIATE								= 11'b01000110000,
							XOR_HALFWORD_IMMEDIATE	  						= 11'b01000101000,
							XOR_WORD_IMMEDIATE		  						= 11'b01000100000,
							FLOATING_ADD									= 11'b01011000100,
							FLOATING_SUBTRACT								= 11'b01011000101,
							FLOATING_MULTIPLY         						= 11'b01011000110,
							FLOATING_MULTIPLY_AND_ADD 						= 11'b11100000000,
							FLOATING_MULTIPLY_AND_SUBTRACT  				= 11'b11110000000,
							EQUIVALENT										= 11'b01001001001,
							SHIFT_LEFT_HALFWORD								= 11'b00001011111,
							SHIFT_LEFT_HALFWORD_IMMEDIATE   				= 11'b00001111111,
							SHIFT_LEFT_WORD									= 11'b00001011011,
							SHIFT_LEFT_WORD_IMMEDIATE						= 11'b00001111011,
							ROTATE_HALFWORD									= 11'b00001011100,
							ROTATE_HALFWORD_IMMEDIATE						= 11'b00001111100,
							ROTATE_WORD										= 11'b00001011000,
							ROTATE_WORD_IMMEDIATE							= 11'b00001111000,
							ROTATE_AND_MASK_HALFWORD						= 11'b00001011101,
							ROTATE_AND_MASK_HALFWORD_IMMEDIATE 				= 11'b00001111101,
							COUNT_ONES_IN_BYTES				   				= 11'b01010110100,
							AVERAGE_BYTES					   				= 11'b00011010011,
							ABSOLUTE_DIFFERENCE_OF_BYTES	  				= 11'b00001010011,
							SUM_BYTES_INTO_HALFWORDS		   				= 11'b01001010011,
							COMPARE_EQUAL_HALFWORD			   				= 11'b01111001000,
							COMPARE_EQUAL_HALFWORD_IMMEDIATE   				= 11'b01111101000,
							COMPARE_EQUAL_WORD				   				= 11'b01111000000,
							COMPARE_EQUAL_WORD_IMMEDIATE	   				= 11'b01111100000,
							COMPARE_GREATER_THAN_HALFWORD      				= 11'b01001001000,
							COMPARE_GREATER_THAN_HALFWORD_IMMEDIATE			= 11'b01001101000,
							COMPARE_GREATER_THAN_WORD						= 11'b01001000000,
							COMPARE_GREATER_THAN_WORD_IMMEDIATE	    		= 11'b01001100000,
							COMPARE_LOGICAL_GREATER_THAN_WORD				= 11'b01011000000,
							COMPARE_LOGICAL_GREATER_THAN_WORD_IMMEDIATE		= 11'b01011100000,
							COMPARE_LOGICAL_GREATER_THAN_HALFWORD		    = 11'b01011001000,
							COMPARE_LOGICAL_GREATER_THAN_HALFWORD_IMMEDIATE = 11'b01011101000,
							CARRY_GENERATE									= 11'b00011000010,
							ADD_EXTENDED									= 11'b01101000000,
							BORROW_GENERATE									= 11'b00001000010,
							SUBTRACT_FROM_EXTENDED							= 11'b01101000001,
							NOP_LOAD										= 11'b00000000001,
							NOP_EXEC 										= 11'b01000000001,
							STOP_AND_SIGNAL									= 11'b00000000000,
							
							LOAD_QUADWORD_DFORM								= 11'b00110100000,
							LOAD_QUADWORD_AFORM 							= 11'b00110000100,
							STORE_QUADWORD_DFORM							= 11'b00100100000,
							STORE_QUADWORD_AFORM							= 11'b00100000100,
							IMMEDIATE_LOAD_HALFWORD							= 11'b01000001100,
							IMMEDIATE_LOAD_WORD								= 11'b01000000100,
							IMMEDIATE_LOAD_ADDRESS							= 11'b01000010000,
							GATHER_BITS_FROM_WORDS							= 11'b00110110000,
							GATHER_BITS_FROM_HALFWORDS						= 11'b00110110001,
							SHUFFLE_BYTES			  						= 11'b10110000000,
							SHIFT_LEFT_QUADWORD_BY_BITS						= 11'b00111011011,
							SHIFT_LEFT_QUADWORD_BY_BITS_IMMEDIATE			= 11'b00111111011,
							SHIFT_LEFT_QUADWORD_BY_BYTES					= 11'b00111011111,
							SHIFT_LEFT_QUADWORD_BY_BYTES_IMMEDIATE			= 11'b00111111111,
							ROTATE_QUADWORD_BY_BYTES						= 11'b00111011100,
							ROTATE_QUADWORD_BY_BYTES_IMMEDIATE				= 11'b00111111100,
							BRANCH_RELATIVE									= 11'b00110010000,
							BRANCH_ABSOLUTE									= 11'b00110000000,
							BRANCH_IF_NOT_ZERO_WORD							= 11'b00100001000,
							BRANCH_IF_ZERO_WORD								= 11'b00100000000,
							BRANCH_IF_NOT_ZERO_HALFWORD						= 11'b00100011000,
							BRANCH_IF_ZERO_HALFWORD							= 11'b00100010000,
							BRANCH_RELATIVE_AND_SET_LINK					= 11'b00110011000,
							BRANCH_ABSOLUTE_AND_SET_LINK					= 11'b00110001000
							} opcode;
							
		parameter LS_SIZE = 320000;
							
endpackage
							
							